localparam [63 : 0] C [0 : 23] = {64'h3BF5080AC8BA94B1,
                                  64'hC1D1659C1BBD92F6,
                                  64'h60E8B2CE0DDEC97B,
                                  64'hEC5FB8FE790FBC13,
                                  64'hAA043DE6436706A7,
                                  64'h8929FF6A5E535BFD,
                                  64'h98BF1E2C50C97550,
                                  64'h4C5F8F162864BAA8,
                                  64'h262FC78B14325D54,
                                  64'h1317E3C58A192EAA,
                                  64'h098BF1E2C50C9755,
                                  64'hD8EE19681D669304,
                                  64'h6C770CB40EB34982,
                                  64'h363B865A0759A4C1,
                                  64'hC73622B47C4C0ACE,
                                  64'h639B115A3E260567,
                                  64'hEDE6693460F3DA1D,
                                  64'hAAD8D5034F9935A0,
                                  64'h556C6A81A7CC9AD0,
                                  64'h2AB63540D3E64D68,
                                  64'h155B1AA069F326B4,
                                  64'h0AAD8D5034F9935A,
                                  64'h0556C6A81A7CC9AD,
                                  64'hDE8082CD72DEBC78};

localparam [5 : 0] M1 [0 : 7] = {6'd8,  6'd56, 6'd8,  6'd56, 6'd8,  6'd56, 6'd8,  6'd56};
localparam [5 : 0] N1 [0 : 7] = {6'd53, 6'd51, 6'd37, 6'd3,  6'd21, 6'd19, 6'd5,  6'd35};
localparam [5 : 0] M2 [0 : 7] = {6'd14, 6'd34, 6'd46, 6'd2,  6'd14, 6'd34, 6'd46, 6'd2};
localparam [5 : 0] N2 [0 : 7] = {6'd1,  6'd7,  6'd49, 6'd23, 6'd33, 6'd39, 6'd17, 6'd55};
