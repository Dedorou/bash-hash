package tb_pkg;

import bash_hash_params_pkg::*;

// bash-s
localparam logic [SLEN-1:0] bash_s_i [0:2] = {64'hB194BAC80A08F53B, 64'hE12BDC1AE28257EC, 64'hE9DEE72C8F0C0FA6};
localparam logic [SLEN-1:0] bash_s_o [0:2] = {64'h479E76129979DC5F, 64'h0F2B2C93ED128EDD, 64'h41009B1B112DFEF3};

localparam logic [5:0] bash_s_param [0:3] = {6'd8, 6'd53, 6'd14, 6'd1};

localparam logic [SLEN-1:0] bash_f_i [0:23] = {64'hB194BAC80A08F53B, 64'h366D008E584A5DE4, 64'h8504FA9D1BB6C7AC, 64'h252E72C202FDCE0D,
                                               64'h5BE3D61217B96181, 64'hFE6786AD716B890B, 64'h5CB0C0FF33C356B8, 64'h35C405AED8E07F99,
                                               64'hE12BDC1AE28257EC, 64'h703FCCF095EE8DF1, 64'hC1AB76389FE678CA, 64'hF7C6F860D5BB9C4F,
                                               64'hF33C657B637C306A, 64'hDD4EA7799EB23D31, 64'h3E98B56E27D3BCCF, 64'h591E181F4C5AB793,
                                               64'hE9DEE72C8F0C0FA6, 64'h2DDB49F46F739647, 64'h06075316ED247A37, 64'h39CBA38303A98BF6,
                                               64'h92BD9B1CE5D14101, 64'h5445FBC95E4D0EF2, 64'h682080AA227D642F, 64'h2687F93490405511};

localparam logic [SLEN-1:0] bash_f_o [0:23] = {64'h8FE727775EA7F140, 64'hB95BB6A200CBB28C, 64'h7F0809C0C0BC68B7, 64'hDC5AEDC841BD94E4,
                                               64'h03630C301FC255DF, 64'h5B67DB53EF65E376, 64'hE8A4D797A6172F22, 64'h71BA48093173D329,
                                               64'hC3502AC946767326, 64'hA2891971392D3F70, 64'h89959F5D61621238, 64'h655975E00E2132A0,
                                               64'hD5018CEEDB17731C, 64'hCD88FC50151D37C0, 64'hD4A3359506AEDC2E, 64'h6109511E7703AFBB,
                                               64'h014642348D8568AA, 64'h1A5D9868C4C7E6DF, 64'hA756B1690C7C2608, 64'hA2DC136F5997AB8F,
                                               64'hBB3F4D9F033C87CA, 64'h6070E117F099C409, 64'h4972ACD9D976214B, 64'h7CED8E3F8B6E058E};

endpackage : tb_pkg

